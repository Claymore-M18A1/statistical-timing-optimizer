module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire net118;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire _426_;
 wire _427_;
 wire _428_;
 wire _429_;
 wire _430_;
 wire _431_;
 wire _432_;
 wire _433_;
 wire _434_;
 wire _435_;
 wire _436_;
 wire _437_;
 wire _438_;
 wire _439_;
 wire _440_;
 wire _441_;
 wire _442_;
 wire _443_;
 wire _444_;
 wire _445_;
 wire _446_;
 wire _447_;
 wire _448_;
 wire _449_;
 wire _450_;
 wire _451_;
 wire _452_;
 wire _453_;
 wire _454_;
 wire _455_;
 wire _456_;
 wire _457_;
 wire _458_;
 wire _459_;
 wire _460_;
 wire _461_;
 wire _462_;
 wire _463_;
 wire _464_;
 wire _465_;
 wire _466_;
 wire _467_;
 wire _468_;
 wire _469_;
 wire _470_;
 wire _471_;
 wire _472_;
 wire _473_;
 wire _474_;
 wire _475_;
 wire _476_;
 wire _477_;
 wire _478_;
 wire _479_;
 wire _480_;
 wire _481_;
 wire _482_;
 wire _483_;
 wire _484_;
 wire _485_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net72;
 wire net73;
 wire net74;
 wire net80;
 wire net81;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net75;
 wire net76;
 wire net77;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net94;
 wire net97;

 INV_X2 _486_ (.A(\dpath.a_lt_b$in1[11] ),
    .ZN(_036_));
 INV_X2 _487_ (.A(\dpath.a_lt_b$in1[10] ),
    .ZN(_037_));
 INV_X2 _488_ (.A(\dpath.a_lt_b$in1[9] ),
    .ZN(_038_));
 INV_X4 _489_ (.A(\dpath.a_lt_b$in1[8] ),
    .ZN(_039_));
 NAND4_X2 _490_ (.A1(_036_),
    .A2(net73),
    .A3(net89),
    .A4(net85),
    .ZN(_040_));
 INV_X1 _491_ (.A(\dpath.a_lt_b$in1[15] ),
    .ZN(_041_));
 INV_X1 _492_ (.A(\dpath.a_lt_b$in1[14] ),
    .ZN(_042_));
 INV_X1 _493_ (.A(\dpath.a_lt_b$in1[13] ),
    .ZN(_043_));
 INV_X2 _494_ (.A(\dpath.a_lt_b$in1[12] ),
    .ZN(_044_));
 NAND4_X2 _495_ (.A1(_041_),
    .A2(_042_),
    .A3(_043_),
    .A4(net68),
    .ZN(_045_));
 INV_X2 _496_ (.A(\dpath.a_lt_b$in1[3] ),
    .ZN(_046_));
 INV_X2 _497_ (.A(\dpath.a_lt_b$in1[2] ),
    .ZN(_047_));
 INV_X2 _498_ (.A(\dpath.a_lt_b$in1[1] ),
    .ZN(_048_));
 INV_X2 _499_ (.A(\dpath.a_lt_b$in1[0] ),
    .ZN(_049_));
 NAND4_X1 _500_ (.A1(_046_),
    .A2(_047_),
    .A3(_048_),
    .A4(_049_),
    .ZN(_050_));
 INV_X2 _501_ (.A(\dpath.a_lt_b$in1[7] ),
    .ZN(_051_));
 INV_X2 _502_ (.A(\dpath.a_lt_b$in1[6] ),
    .ZN(_052_));
 INV_X2 _503_ (.A(\dpath.a_lt_b$in1[5] ),
    .ZN(_053_));
 INV_X2 _504_ (.A(\dpath.a_lt_b$in1[4] ),
    .ZN(_054_));
 NAND4_X2 _505_ (.A1(_051_),
    .A2(net123),
    .A3(net103),
    .A4(net101),
    .ZN(_055_));
 NOR4_X1 _506_ (.A1(_040_),
    .A2(_045_),
    .A3(_050_),
    .A4(_055_),
    .ZN(_056_));
 BUF_X4 _507_ (.A(\ctrl.state.out[2] ),
    .Z(_057_));
 INV_X2 _508_ (.A(_057_),
    .ZN(_058_));
 OR2_X1 _509_ (.A1(_058_),
    .A2(net34),
    .ZN(_059_));
 BUF_X4 _510_ (.A(net36),
    .Z(_060_));
 BUF_X4 _511_ (.A(_060_),
    .Z(_061_));
 BUF_X4 _512_ (.A(_061_),
    .Z(_062_));
 NAND2_X1 _513_ (.A1(_062_),
    .A2(net33),
    .ZN(_063_));
 OAI22_X1 _514_ (.A1(_056_),
    .A2(_059_),
    .B1(net34),
    .B2(_063_),
    .ZN(_002_));
 BUF_X2 _515_ (.A(_003_),
    .Z(_064_));
 AND3_X2 _516_ (.A1(_058_),
    .A2(\ctrl.state.out[1] ),
    .A3(_064_),
    .ZN(net53));
 AOI21_X2 _517_ (.A(net34),
    .B1(net53),
    .B2(net35),
    .ZN(_065_));
 BUF_X4 _518_ (.A(_060_),
    .Z(_066_));
 BUF_X2 _519_ (.A(_066_),
    .Z(_067_));
 INV_X1 _520_ (.A(_067_),
    .ZN(_068_));
 OAI21_X2 _521_ (.A(_065_),
    .B1(_068_),
    .B2(net33),
    .ZN(_000_));
 NAND2_X1 _522_ (.A1(_065_),
    .A2(\ctrl.state.out[1] ),
    .ZN(_069_));
 INV_X2 _523_ (.A(_056_),
    .ZN(_070_));
 OAI21_X1 _524_ (.A(_069_),
    .B1(_070_),
    .B2(_059_),
    .ZN(_001_));
 XNOR2_X1 _525_ (.A(_049_),
    .B(\dpath.a_lt_b$in0[0] ),
    .ZN(net37));
 BUF_X2 rebuffer65 (.A(_081_),
    .Z(net118));
 NAND2_X2 _527_ (.A1(_048_),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_072_));
 NOR2_X2 _528_ (.A1(_049_),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_073_));
 NOR2_X2 _529_ (.A1(_048_),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_074_));
 OAI21_X2 _530_ (.A(_072_),
    .B1(_073_),
    .B2(_074_),
    .ZN(_075_));
 NAND2_X2 _531_ (.A1(_046_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_076_));
 INV_X2 _532_ (.A(\dpath.a_lt_b$in0[3] ),
    .ZN(_077_));
 NAND2_X4 _533_ (.A1(_077_),
    .A2(net119),
    .ZN(_078_));
 NAND2_X4 _534_ (.A1(_078_),
    .A2(_076_),
    .ZN(_079_));
 NAND2_X2 _535_ (.A1(_047_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_080_));
 INV_X2 _536_ (.A(\dpath.a_lt_b$in0[2] ),
    .ZN(_081_));
 NAND2_X4 _537_ (.A1(_081_),
    .A2(net117),
    .ZN(_082_));
 NAND2_X4 _538_ (.A1(_082_),
    .A2(_080_),
    .ZN(_083_));
 NOR2_X2 _539_ (.A1(_083_),
    .A2(_079_),
    .ZN(_084_));
 NAND2_X4 _540_ (.A1(_075_),
    .A2(_084_),
    .ZN(_085_));
 NOR2_X2 _541_ (.A1(_046_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_086_));
 OAI21_X2 _542_ (.A(_076_),
    .B1(_086_),
    .B2(_080_),
    .ZN(_087_));
 INV_X1 _543_ (.A(_087_),
    .ZN(_088_));
 NAND2_X4 _544_ (.A1(_085_),
    .A2(_088_),
    .ZN(_089_));
 INV_X1 _545_ (.A(\dpath.a_lt_b$in0[7] ),
    .ZN(_090_));
 NAND2_X2 _546_ (.A1(_090_),
    .A2(\dpath.a_lt_b$in1[7] ),
    .ZN(_091_));
 NAND2_X4 _547_ (.A1(_051_),
    .A2(net75),
    .ZN(_092_));
 NAND2_X4 _548_ (.A1(_091_),
    .A2(_092_),
    .ZN(_093_));
 NAND2_X4 _549_ (.A1(_052_),
    .A2(\dpath.a_lt_b$in0[6] ),
    .ZN(_094_));
 INV_X2 _550_ (.A(\dpath.a_lt_b$in0[6] ),
    .ZN(_095_));
 NAND2_X4 _551_ (.A1(_095_),
    .A2(\dpath.a_lt_b$in1[6] ),
    .ZN(_096_));
 NAND2_X4 _552_ (.A1(_094_),
    .A2(_096_),
    .ZN(_097_));
 NOR2_X4 _553_ (.A1(_097_),
    .A2(_093_),
    .ZN(_098_));
 NAND2_X4 _554_ (.A1(_053_),
    .A2(\dpath.a_lt_b$in0[5] ),
    .ZN(_099_));
 INV_X2 _555_ (.A(\dpath.a_lt_b$in0[5] ),
    .ZN(_100_));
 NAND2_X4 _556_ (.A1(_100_),
    .A2(\dpath.a_lt_b$in1[5] ),
    .ZN(_101_));
 NAND2_X4 _557_ (.A1(_101_),
    .A2(_099_),
    .ZN(_102_));
 NAND2_X4 _558_ (.A1(net62),
    .A2(_054_),
    .ZN(_103_));
 INV_X2 _559_ (.A(\dpath.a_lt_b$in0[4] ),
    .ZN(_104_));
 NAND2_X2 _560_ (.A1(_104_),
    .A2(net77),
    .ZN(_105_));
 NAND2_X2 _561_ (.A1(_103_),
    .A2(_105_),
    .ZN(_106_));
 NOR2_X4 _562_ (.A1(_102_),
    .A2(_106_),
    .ZN(_107_));
 AND2_X4 _563_ (.A1(_098_),
    .A2(_107_),
    .ZN(_108_));
 NAND2_X4 _564_ (.A1(net116),
    .A2(_108_),
    .ZN(_109_));
 NAND2_X2 _565_ (.A1(_092_),
    .A2(_094_),
    .ZN(_110_));
 NAND2_X2 _566_ (.A1(_110_),
    .A2(_091_),
    .ZN(_111_));
 INV_X2 _567_ (.A(_111_),
    .ZN(_112_));
 INV_X1 _568_ (.A(_099_),
    .ZN(_113_));
 NOR2_X2 _569_ (.A1(_104_),
    .A2(\dpath.a_lt_b$in1[4] ),
    .ZN(_114_));
 OAI21_X4 _570_ (.A(net57),
    .B1(_113_),
    .B2(_114_),
    .ZN(_115_));
 INV_X1 _571_ (.A(_115_),
    .ZN(_116_));
 AOI21_X2 _572_ (.A(_112_),
    .B1(_116_),
    .B2(_098_),
    .ZN(_117_));
 NAND2_X2 _573_ (.A1(_109_),
    .A2(_117_),
    .ZN(_118_));
 INV_X1 _574_ (.A(\dpath.a_lt_b$in0[13] ),
    .ZN(_119_));
 NOR2_X2 _575_ (.A1(_119_),
    .A2(\dpath.a_lt_b$in1[13] ),
    .ZN(_120_));
 INV_X1 _576_ (.A(_120_),
    .ZN(_121_));
 NAND2_X2 _577_ (.A1(_119_),
    .A2(\dpath.a_lt_b$in1[13] ),
    .ZN(_122_));
 NAND2_X2 _578_ (.A1(_121_),
    .A2(_122_),
    .ZN(_123_));
 INV_X2 _579_ (.A(_123_),
    .ZN(_124_));
 INV_X2 _580_ (.A(\dpath.a_lt_b$in0[12] ),
    .ZN(_125_));
 NOR2_X4 _581_ (.A1(_125_),
    .A2(\dpath.a_lt_b$in1[12] ),
    .ZN(_126_));
 NOR2_X4 _582_ (.A1(_044_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_127_));
 NOR2_X4 _583_ (.A1(_126_),
    .A2(_127_),
    .ZN(_128_));
 NAND2_X1 _584_ (.A1(_124_),
    .A2(_128_),
    .ZN(_129_));
 NAND2_X2 _585_ (.A1(_042_),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_130_));
 INV_X2 _586_ (.A(\dpath.a_lt_b$in0[14] ),
    .ZN(_131_));
 NAND2_X2 _587_ (.A1(_131_),
    .A2(\dpath.a_lt_b$in1[14] ),
    .ZN(_132_));
 NAND2_X2 _588_ (.A1(_130_),
    .A2(_132_),
    .ZN(_133_));
 INV_X1 _589_ (.A(_133_),
    .ZN(_134_));
 XNOR2_X1 _590_ (.A(\dpath.a_lt_b$in1[15] ),
    .B(\dpath.a_lt_b$in0[15] ),
    .ZN(_135_));
 NAND2_X2 _591_ (.A1(_134_),
    .A2(_135_),
    .ZN(_136_));
 NOR2_X2 _592_ (.A1(_129_),
    .A2(_136_),
    .ZN(_137_));
 NAND2_X4 _593_ (.A1(_036_),
    .A2(net81),
    .ZN(_138_));
 INV_X2 _594_ (.A(\dpath.a_lt_b$in0[11] ),
    .ZN(_139_));
 NAND2_X2 _595_ (.A1(_139_),
    .A2(\dpath.a_lt_b$in1[11] ),
    .ZN(_140_));
 NAND2_X2 _596_ (.A1(_138_),
    .A2(_140_),
    .ZN(_141_));
 NAND2_X4 _597_ (.A1(_037_),
    .A2(net64),
    .ZN(_142_));
 INV_X2 _598_ (.A(\dpath.a_lt_b$in0[10] ),
    .ZN(_143_));
 NAND2_X2 _599_ (.A1(_143_),
    .A2(\dpath.a_lt_b$in1[10] ),
    .ZN(_144_));
 NAND2_X4 _600_ (.A1(_142_),
    .A2(_144_),
    .ZN(_145_));
 NOR2_X4 _601_ (.A1(_141_),
    .A2(_145_),
    .ZN(_146_));
 INV_X2 _602_ (.A(_146_),
    .ZN(_147_));
 NAND2_X4 _603_ (.A1(_038_),
    .A2(net72),
    .ZN(_148_));
 INV_X2 _604_ (.A(\dpath.a_lt_b$in0[9] ),
    .ZN(_149_));
 NAND2_X2 _605_ (.A1(_149_),
    .A2(\dpath.a_lt_b$in1[9] ),
    .ZN(_150_));
 NAND2_X2 _606_ (.A1(_148_),
    .A2(_150_),
    .ZN(_151_));
 INV_X4 _607_ (.A(_151_),
    .ZN(_152_));
 NAND2_X2 _608_ (.A1(_039_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_153_));
 INV_X2 _609_ (.A(\dpath.a_lt_b$in0[8] ),
    .ZN(_154_));
 NAND2_X4 _610_ (.A1(_154_),
    .A2(\dpath.a_lt_b$in1[8] ),
    .ZN(_155_));
 NAND2_X4 _611_ (.A1(_153_),
    .A2(_155_),
    .ZN(_156_));
 INV_X4 _612_ (.A(_156_),
    .ZN(_157_));
 NAND2_X2 _613_ (.A1(_152_),
    .A2(_157_),
    .ZN(_158_));
 NOR2_X2 _614_ (.A1(_158_),
    .A2(_147_),
    .ZN(_159_));
 AND2_X2 _615_ (.A1(_137_),
    .A2(net80),
    .ZN(_160_));
 NAND2_X4 _616_ (.A1(net114),
    .A2(_160_),
    .ZN(_161_));
 NAND2_X1 _617_ (.A1(_148_),
    .A2(_153_),
    .ZN(_162_));
 NAND2_X1 _618_ (.A1(_162_),
    .A2(_150_),
    .ZN(_163_));
 INV_X1 _619_ (.A(_163_),
    .ZN(_164_));
 NAND2_X2 _620_ (.A1(_146_),
    .A2(_164_),
    .ZN(_165_));
 INV_X2 _621_ (.A(_138_),
    .ZN(_166_));
 INV_X1 _622_ (.A(_142_),
    .ZN(_167_));
 OAI21_X1 _623_ (.A(_140_),
    .B1(_166_),
    .B2(_167_),
    .ZN(_168_));
 NAND2_X2 _624_ (.A1(_165_),
    .A2(_168_),
    .ZN(_169_));
 NAND2_X1 _625_ (.A1(_169_),
    .A2(_137_),
    .ZN(_170_));
 OAI21_X1 _626_ (.A(_122_),
    .B1(_120_),
    .B2(_126_),
    .ZN(_171_));
 NOR2_X1 _627_ (.A1(_171_),
    .A2(_136_),
    .ZN(_172_));
 NAND2_X1 _628_ (.A1(_041_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_173_));
 INV_X1 _629_ (.A(_135_),
    .ZN(_174_));
 OAI21_X2 _630_ (.A(_173_),
    .B1(_174_),
    .B2(_130_),
    .ZN(_175_));
 NOR2_X1 _631_ (.A1(_172_),
    .A2(_175_),
    .ZN(_176_));
 NAND2_X1 _632_ (.A1(_170_),
    .A2(_176_),
    .ZN(_177_));
 INV_X4 _633_ (.A(_177_),
    .ZN(_178_));
 NAND2_X4 _634_ (.A1(_161_),
    .A2(_178_),
    .ZN(_179_));
 NAND2_X2 _635_ (.A1(_057_),
    .A2(_003_),
    .ZN(_180_));
 INV_X4 _636_ (.A(_180_),
    .ZN(_181_));
 NAND3_X1 _637_ (.A1(_179_),
    .A2(net37),
    .A3(_181_),
    .ZN(_182_));
 NAND4_X2 _638_ (.A1(_161_),
    .A2(_057_),
    .A3(_064_),
    .A4(_178_),
    .ZN(_183_));
 OAI21_X1 _639_ (.A(_182_),
    .B1(_183_),
    .B2(_049_),
    .ZN(_184_));
 NOR2_X2 _640_ (.A1(_058_),
    .A2(_060_),
    .ZN(_185_));
 BUF_X4 _641_ (.A(_185_),
    .Z(_186_));
 NAND2_X1 _642_ (.A1(_184_),
    .A2(_186_),
    .ZN(_187_));
 NOR2_X2 _643_ (.A1(_060_),
    .A2(_057_),
    .ZN(_188_));
 BUF_X2 _644_ (.A(_188_),
    .Z(_189_));
 AND2_X1 _645_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_190_));
 AOI21_X1 _646_ (.A(_190_),
    .B1(_067_),
    .B2(net8),
    .ZN(_191_));
 NAND2_X1 _647_ (.A1(_187_),
    .A2(_191_),
    .ZN(_004_));
 NAND3_X2 _648_ (.A1(_161_),
    .A2(_057_),
    .A3(_178_),
    .ZN(_192_));
 INV_X2 _649_ (.A(_192_),
    .ZN(_193_));
 NAND3_X1 _650_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[10] ),
    .A3(_064_),
    .ZN(_194_));
 NAND2_X4 _651_ (.A1(_107_),
    .A2(_087_),
    .ZN(_195_));
 NAND2_X4 _652_ (.A1(_195_),
    .A2(_115_),
    .ZN(_196_));
 INV_X4 _653_ (.A(_196_),
    .ZN(_197_));
 NAND3_X2 _654_ (.A1(_075_),
    .A2(_084_),
    .A3(_107_),
    .ZN(_198_));
 NAND2_X4 _655_ (.A1(_197_),
    .A2(_198_),
    .ZN(_199_));
 NAND3_X2 _656_ (.A1(_098_),
    .A2(_152_),
    .A3(net60),
    .ZN(_200_));
 INV_X2 _657_ (.A(_200_),
    .ZN(_201_));
 NAND2_X4 _658_ (.A1(_199_),
    .A2(_201_),
    .ZN(_202_));
 OAI21_X2 _659_ (.A(_163_),
    .B1(_158_),
    .B2(_111_),
    .ZN(_203_));
 INV_X2 _660_ (.A(_203_),
    .ZN(_204_));
 NAND2_X2 _661_ (.A1(_204_),
    .A2(_202_),
    .ZN(_205_));
 XNOR2_X2 _662_ (.A(_145_),
    .B(_205_),
    .ZN(net38));
 AOI21_X4 _663_ (.A(_180_),
    .B1(_161_),
    .B2(_178_),
    .ZN(_206_));
 NAND2_X1 _664_ (.A1(net76),
    .A2(_206_),
    .ZN(_207_));
 NAND2_X1 _665_ (.A1(_194_),
    .A2(_207_),
    .ZN(_208_));
 NAND2_X1 _666_ (.A1(_208_),
    .A2(_186_),
    .ZN(_209_));
 AND2_X2 _667_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[10] ),
    .ZN(_210_));
 AOI21_X1 _668_ (.A(_210_),
    .B1(_067_),
    .B2(net19),
    .ZN(_211_));
 NAND2_X1 _669_ (.A1(_209_),
    .A2(_211_),
    .ZN(_005_));
 NAND3_X2 _670_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[11] ),
    .A3(_064_),
    .ZN(_212_));
 INV_X2 _671_ (.A(_083_),
    .ZN(_213_));
 XNOR2_X2 _672_ (.A(\dpath.a_lt_b$in1[1] ),
    .B(\dpath.a_lt_b$in0[1] ),
    .ZN(_214_));
 INV_X2 _673_ (.A(_073_),
    .ZN(_215_));
 NAND3_X4 _674_ (.A1(_214_),
    .A2(_213_),
    .A3(_215_),
    .ZN(_216_));
 NOR2_X1 _675_ (.A1(_047_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_217_));
 OAI21_X2 _676_ (.A(_080_),
    .B1(_217_),
    .B2(_072_),
    .ZN(_218_));
 INV_X1 _677_ (.A(_218_),
    .ZN(_219_));
 NAND2_X2 _678_ (.A1(_216_),
    .A2(_219_),
    .ZN(_220_));
 NOR2_X4 _679_ (.A1(_106_),
    .A2(_079_),
    .ZN(_221_));
 INV_X2 _680_ (.A(_221_),
    .ZN(_222_));
 NOR2_X2 _681_ (.A1(_102_),
    .A2(_097_),
    .ZN(_223_));
 INV_X4 _682_ (.A(_223_),
    .ZN(_224_));
 NOR2_X2 _683_ (.A1(_224_),
    .A2(_222_),
    .ZN(_225_));
 NAND2_X4 _684_ (.A1(_225_),
    .A2(_220_),
    .ZN(_226_));
 NAND2_X1 _685_ (.A1(_094_),
    .A2(_099_),
    .ZN(_227_));
 NAND2_X2 _686_ (.A1(_227_),
    .A2(_096_),
    .ZN(_228_));
 INV_X2 _687_ (.A(_228_),
    .ZN(_229_));
 INV_X2 _688_ (.A(_076_),
    .ZN(_230_));
 OAI21_X2 _689_ (.A(_105_),
    .B1(_230_),
    .B2(_114_),
    .ZN(_231_));
 INV_X2 _690_ (.A(_231_),
    .ZN(_232_));
 AOI21_X4 _691_ (.A(_229_),
    .B1(_232_),
    .B2(net61),
    .ZN(_233_));
 NAND2_X2 _692_ (.A1(_226_),
    .A2(_233_),
    .ZN(_234_));
 INV_X1 _693_ (.A(_145_),
    .ZN(_235_));
 NAND2_X2 _694_ (.A1(_235_),
    .A2(_152_),
    .ZN(_236_));
 INV_X1 _695_ (.A(_236_),
    .ZN(_237_));
 INV_X4 _696_ (.A(_093_),
    .ZN(_238_));
 NAND2_X4 _697_ (.A1(_238_),
    .A2(_157_),
    .ZN(_239_));
 INV_X2 _698_ (.A(_239_),
    .ZN(_240_));
 NAND2_X2 _699_ (.A1(_237_),
    .A2(_240_),
    .ZN(_241_));
 INV_X2 _700_ (.A(_241_),
    .ZN(_242_));
 NAND2_X1 _701_ (.A1(_234_),
    .A2(_242_),
    .ZN(_243_));
 INV_X2 _702_ (.A(_148_),
    .ZN(_244_));
 OAI21_X2 _703_ (.A(net74),
    .B1(_167_),
    .B2(_244_),
    .ZN(_245_));
 NAND2_X2 _704_ (.A1(_092_),
    .A2(_153_),
    .ZN(_246_));
 NAND2_X1 _705_ (.A1(_246_),
    .A2(net84),
    .ZN(_247_));
 OAI21_X1 _706_ (.A(_245_),
    .B1(_236_),
    .B2(_247_),
    .ZN(_248_));
 INV_X1 _707_ (.A(_248_),
    .ZN(_249_));
 NAND2_X2 _708_ (.A1(_243_),
    .A2(_249_),
    .ZN(_250_));
 NAND2_X1 _709_ (.A1(_250_),
    .A2(_141_),
    .ZN(_251_));
 INV_X1 _710_ (.A(_141_),
    .ZN(_252_));
 NAND3_X2 _711_ (.A1(_243_),
    .A2(_252_),
    .A3(_249_),
    .ZN(_253_));
 NAND2_X2 _712_ (.A1(_251_),
    .A2(_253_),
    .ZN(net39));
 NAND2_X2 _713_ (.A1(net39),
    .A2(_206_),
    .ZN(_254_));
 NAND2_X1 _714_ (.A1(_212_),
    .A2(_254_),
    .ZN(_255_));
 NAND2_X1 _715_ (.A1(_255_),
    .A2(_186_),
    .ZN(_256_));
 AND2_X2 _716_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_257_));
 AOI21_X2 _717_ (.A(_257_),
    .B1(_067_),
    .B2(net20),
    .ZN(_258_));
 NAND2_X1 _718_ (.A1(_256_),
    .A2(_258_),
    .ZN(_006_));
 NAND3_X1 _719_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[12] ),
    .A3(_064_),
    .ZN(_259_));
 INV_X1 _720_ (.A(_098_),
    .ZN(_260_));
 OAI21_X2 _721_ (.A(_111_),
    .B1(_260_),
    .B2(_115_),
    .ZN(_261_));
 NAND2_X1 _722_ (.A1(_261_),
    .A2(_159_),
    .ZN(_262_));
 INV_X1 _723_ (.A(_169_),
    .ZN(_263_));
 NAND2_X2 _724_ (.A1(_262_),
    .A2(_263_),
    .ZN(_264_));
 NAND2_X4 _725_ (.A1(_108_),
    .A2(_159_),
    .ZN(_265_));
 INV_X1 _726_ (.A(_089_),
    .ZN(_266_));
 NOR2_X4 _727_ (.A1(_266_),
    .A2(_265_),
    .ZN(_267_));
 NOR2_X2 _728_ (.A1(_267_),
    .A2(_264_),
    .ZN(_268_));
 NAND2_X1 _729_ (.A1(net55),
    .A2(_268_),
    .ZN(_269_));
 INV_X4 _730_ (.A(_128_),
    .ZN(_270_));
 OAI21_X2 _731_ (.A(_270_),
    .B1(_264_),
    .B2(_267_),
    .ZN(_271_));
 NAND2_X2 _732_ (.A1(_269_),
    .A2(_271_),
    .ZN(net40));
 NAND2_X2 _733_ (.A1(net94),
    .A2(_206_),
    .ZN(_272_));
 NAND2_X1 _734_ (.A1(_259_),
    .A2(_272_),
    .ZN(_273_));
 NAND2_X1 _735_ (.A1(_273_),
    .A2(_186_),
    .ZN(_274_));
 AND2_X2 _736_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_275_));
 AOI21_X2 _737_ (.A(_275_),
    .B1(_067_),
    .B2(net21),
    .ZN(_276_));
 NAND2_X1 _738_ (.A1(_274_),
    .A2(_276_),
    .ZN(_007_));
 NAND3_X1 _739_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[13] ),
    .A3(_064_),
    .ZN(_277_));
 NOR2_X4 _740_ (.A1(_270_),
    .A2(_141_),
    .ZN(_278_));
 INV_X1 _741_ (.A(_278_),
    .ZN(_279_));
 NOR2_X2 _742_ (.A1(_236_),
    .A2(_279_),
    .ZN(_280_));
 NOR2_X4 _743_ (.A1(_224_),
    .A2(_239_),
    .ZN(_281_));
 AND2_X2 _744_ (.A1(_280_),
    .A2(_281_),
    .ZN(_282_));
 NAND2_X2 _745_ (.A1(_220_),
    .A2(net65),
    .ZN(_283_));
 NAND2_X2 _746_ (.A1(_283_),
    .A2(_231_),
    .ZN(_284_));
 NAND2_X2 _747_ (.A1(_282_),
    .A2(_284_),
    .ZN(_285_));
 OAI21_X1 _748_ (.A(_247_),
    .B1(_239_),
    .B2(_228_),
    .ZN(_286_));
 NAND2_X1 _749_ (.A1(_280_),
    .A2(_286_),
    .ZN(_287_));
 INV_X2 _750_ (.A(_127_),
    .ZN(_288_));
 OAI21_X1 _751_ (.A(_288_),
    .B1(_166_),
    .B2(_126_),
    .ZN(_289_));
 INV_X1 _752_ (.A(_289_),
    .ZN(_290_));
 INV_X1 _753_ (.A(_245_),
    .ZN(_291_));
 AOI21_X2 _754_ (.A(_290_),
    .B1(_291_),
    .B2(_278_),
    .ZN(_292_));
 NAND2_X2 _755_ (.A1(_287_),
    .A2(_292_),
    .ZN(_293_));
 INV_X2 _756_ (.A(_293_),
    .ZN(_294_));
 NAND2_X2 _757_ (.A1(_285_),
    .A2(_294_),
    .ZN(_295_));
 NAND2_X2 _758_ (.A1(_295_),
    .A2(_123_),
    .ZN(_296_));
 NAND3_X1 _759_ (.A1(_285_),
    .A2(_294_),
    .A3(_124_),
    .ZN(_297_));
 NAND2_X2 _760_ (.A1(_296_),
    .A2(_297_),
    .ZN(net41));
 NAND2_X1 _761_ (.A1(net41),
    .A2(_206_),
    .ZN(_298_));
 NAND2_X1 _762_ (.A1(_277_),
    .A2(_298_),
    .ZN(_299_));
 NAND2_X1 _763_ (.A1(_299_),
    .A2(_186_),
    .ZN(_300_));
 AND2_X2 _764_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[13] ),
    .ZN(_301_));
 AOI21_X1 _765_ (.A(_301_),
    .B1(_067_),
    .B2(net22),
    .ZN(_302_));
 NAND2_X1 _766_ (.A1(_300_),
    .A2(_302_),
    .ZN(_008_));
 NAND3_X2 _767_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[14] ),
    .A3(_064_),
    .ZN(_303_));
 NAND3_X2 _768_ (.A1(_146_),
    .A2(_124_),
    .A3(net54),
    .ZN(_304_));
 NOR2_X2 _769_ (.A1(_200_),
    .A2(_304_),
    .ZN(_305_));
 NAND2_X2 _770_ (.A1(_199_),
    .A2(_305_),
    .ZN(_306_));
 INV_X1 _771_ (.A(_306_),
    .ZN(_307_));
 INV_X2 _772_ (.A(_304_),
    .ZN(_308_));
 NAND2_X1 _773_ (.A1(_203_),
    .A2(_308_),
    .ZN(_309_));
 NOR2_X2 _774_ (.A1(_129_),
    .A2(_168_),
    .ZN(_310_));
 INV_X1 _775_ (.A(_171_),
    .ZN(_311_));
 NOR2_X2 _776_ (.A1(_310_),
    .A2(_311_),
    .ZN(_312_));
 NAND2_X2 _777_ (.A1(_309_),
    .A2(_312_),
    .ZN(_313_));
 OAI21_X2 _778_ (.A(_133_),
    .B1(_307_),
    .B2(_313_),
    .ZN(_314_));
 INV_X1 _779_ (.A(_313_),
    .ZN(_315_));
 NAND3_X1 _780_ (.A1(_315_),
    .A2(_306_),
    .A3(_134_),
    .ZN(_316_));
 NAND2_X1 _781_ (.A1(_314_),
    .A2(_316_),
    .ZN(net42));
 NAND2_X2 _782_ (.A1(net42),
    .A2(_206_),
    .ZN(_317_));
 NAND2_X1 _783_ (.A1(_303_),
    .A2(_317_),
    .ZN(_318_));
 NAND2_X2 _784_ (.A1(_318_),
    .A2(_186_),
    .ZN(_319_));
 AND2_X1 _785_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_320_));
 AOI21_X2 _786_ (.A(_320_),
    .B1(_067_),
    .B2(net24),
    .ZN(_321_));
 NAND2_X1 _787_ (.A1(_319_),
    .A2(_321_),
    .ZN(_009_));
 NAND3_X1 _788_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[15] ),
    .A3(_064_),
    .ZN(_322_));
 NOR2_X2 _789_ (.A1(_123_),
    .A2(_133_),
    .ZN(_323_));
 AND2_X2 _790_ (.A1(_278_),
    .A2(_323_),
    .ZN(_324_));
 AND2_X2 _791_ (.A1(_324_),
    .A2(_242_),
    .ZN(_325_));
 NAND2_X2 _792_ (.A1(_234_),
    .A2(_325_),
    .ZN(_326_));
 NAND2_X1 _793_ (.A1(_324_),
    .A2(_248_),
    .ZN(_327_));
 OAI21_X1 _794_ (.A(_130_),
    .B1(_133_),
    .B2(_121_),
    .ZN(_328_));
 AOI21_X1 _795_ (.A(_328_),
    .B1(_290_),
    .B2(_323_),
    .ZN(_329_));
 NAND2_X2 _796_ (.A1(_327_),
    .A2(_329_),
    .ZN(_330_));
 INV_X1 _797_ (.A(_330_),
    .ZN(_331_));
 NAND2_X2 _798_ (.A1(_326_),
    .A2(_331_),
    .ZN(_332_));
 NAND2_X2 _799_ (.A1(_332_),
    .A2(_174_),
    .ZN(_333_));
 NAND3_X1 _800_ (.A1(_326_),
    .A2(_331_),
    .A3(_135_),
    .ZN(_334_));
 NAND2_X2 _801_ (.A1(_333_),
    .A2(_334_),
    .ZN(net43));
 NAND2_X1 _802_ (.A1(net43),
    .A2(_206_),
    .ZN(_335_));
 NAND2_X1 _803_ (.A1(_322_),
    .A2(_335_),
    .ZN(_336_));
 NAND2_X1 _804_ (.A1(_336_),
    .A2(_186_),
    .ZN(_337_));
 AND2_X2 _805_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_338_));
 AOI21_X1 _806_ (.A(_338_),
    .B1(_067_),
    .B2(net25),
    .ZN(_339_));
 NAND2_X2 _807_ (.A1(_337_),
    .A2(_339_),
    .ZN(_010_));
 XNOR2_X1 _808_ (.A(_214_),
    .B(_215_),
    .ZN(_340_));
 INV_X1 _809_ (.A(_340_),
    .ZN(net44));
 NAND3_X1 _810_ (.A1(_179_),
    .A2(_181_),
    .A3(net44),
    .ZN(_341_));
 OAI21_X1 _811_ (.A(_341_),
    .B1(_183_),
    .B2(_048_),
    .ZN(_342_));
 NAND2_X2 _812_ (.A1(_342_),
    .A2(_186_),
    .ZN(_343_));
 AND2_X2 _813_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_344_));
 AOI21_X1 _814_ (.A(_344_),
    .B1(_067_),
    .B2(net9),
    .ZN(_345_));
 NAND2_X1 _815_ (.A1(_343_),
    .A2(_345_),
    .ZN(_011_));
 XNOR2_X1 _816_ (.A(_075_),
    .B(net63),
    .ZN(net45));
 NAND3_X1 _817_ (.A1(_179_),
    .A2(_181_),
    .A3(net45),
    .ZN(_346_));
 OAI21_X1 _818_ (.A(_346_),
    .B1(_183_),
    .B2(_047_),
    .ZN(_347_));
 NAND2_X1 _819_ (.A1(_347_),
    .A2(_186_),
    .ZN(_348_));
 AND2_X2 _820_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_349_));
 AOI21_X1 _821_ (.A(_349_),
    .B1(_067_),
    .B2(net10),
    .ZN(_350_));
 NAND2_X1 _822_ (.A1(_348_),
    .A2(_350_),
    .ZN(_012_));
 XNOR2_X1 _823_ (.A(_220_),
    .B(net120),
    .ZN(net46));
 NAND3_X1 _824_ (.A1(_179_),
    .A2(_181_),
    .A3(net46),
    .ZN(_351_));
 OAI21_X1 _825_ (.A(_351_),
    .B1(_183_),
    .B2(_046_),
    .ZN(_352_));
 NAND2_X2 _826_ (.A1(_352_),
    .A2(_186_),
    .ZN(_353_));
 AND2_X1 _827_ (.A1(_189_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_354_));
 AOI21_X2 _828_ (.A(_354_),
    .B1(_062_),
    .B2(net11),
    .ZN(_355_));
 NAND2_X2 _829_ (.A1(_353_),
    .A2(_355_),
    .ZN(_013_));
 XNOR2_X1 _830_ (.A(net115),
    .B(net70),
    .ZN(net47));
 NAND3_X1 _831_ (.A1(_179_),
    .A2(_181_),
    .A3(net47),
    .ZN(_356_));
 OAI21_X2 _832_ (.A(_356_),
    .B1(_183_),
    .B2(net100),
    .ZN(_357_));
 NAND2_X1 _833_ (.A1(_357_),
    .A2(_185_),
    .ZN(_358_));
 AND2_X1 _834_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[4] ),
    .ZN(_359_));
 AOI21_X1 _835_ (.A(_359_),
    .B1(_062_),
    .B2(net13),
    .ZN(_360_));
 NAND2_X1 _836_ (.A1(_358_),
    .A2(_360_),
    .ZN(_014_));
 NAND2_X1 _837_ (.A1(_284_),
    .A2(_102_),
    .ZN(_361_));
 INV_X1 _838_ (.A(_102_),
    .ZN(_362_));
 NAND3_X1 _839_ (.A1(_283_),
    .A2(_362_),
    .A3(_231_),
    .ZN(_363_));
 NAND2_X1 _840_ (.A1(_361_),
    .A2(_363_),
    .ZN(net48));
 NAND3_X2 _841_ (.A1(_179_),
    .A2(net48),
    .A3(_181_),
    .ZN(_364_));
 OAI21_X1 _842_ (.A(_364_),
    .B1(_183_),
    .B2(net102),
    .ZN(_365_));
 NAND2_X1 _843_ (.A1(_365_),
    .A2(_185_),
    .ZN(_366_));
 AND2_X1 _844_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[5] ),
    .ZN(_367_));
 AOI21_X2 _845_ (.A(_367_),
    .B1(_062_),
    .B2(net14),
    .ZN(_368_));
 NAND2_X1 _846_ (.A1(_366_),
    .A2(_368_),
    .ZN(_015_));
 XNOR2_X2 _847_ (.A(net71),
    .B(_097_),
    .ZN(net49));
 NAND3_X1 _848_ (.A1(_179_),
    .A2(net49),
    .A3(_181_),
    .ZN(_369_));
 OAI21_X1 _849_ (.A(_369_),
    .B1(_183_),
    .B2(_052_),
    .ZN(_370_));
 NAND2_X1 _850_ (.A1(_370_),
    .A2(_185_),
    .ZN(_371_));
 AND2_X1 _851_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[6] ),
    .ZN(_372_));
 AOI21_X2 _852_ (.A(_372_),
    .B1(_062_),
    .B2(net15),
    .ZN(_373_));
 NAND2_X1 _853_ (.A1(_371_),
    .A2(_373_),
    .ZN(_016_));
 NAND2_X4 _854_ (.A1(net58),
    .A2(_093_),
    .ZN(_374_));
 NAND3_X2 _855_ (.A1(net56),
    .A2(net97),
    .A3(_238_),
    .ZN(_375_));
 NAND2_X2 _856_ (.A1(_374_),
    .A2(_375_),
    .ZN(net50));
 NAND3_X2 _857_ (.A1(_179_),
    .A2(net124),
    .A3(_181_),
    .ZN(_376_));
 OAI21_X1 _858_ (.A(_376_),
    .B1(_183_),
    .B2(_051_),
    .ZN(_377_));
 NAND2_X1 _859_ (.A1(_377_),
    .A2(_185_),
    .ZN(_378_));
 AND2_X2 _860_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[7] ),
    .ZN(_379_));
 AOI21_X2 _861_ (.A(_379_),
    .B1(_062_),
    .B2(net16),
    .ZN(_380_));
 NAND2_X1 _862_ (.A1(_378_),
    .A2(_380_),
    .ZN(_017_));
 NAND2_X2 _863_ (.A1(_118_),
    .A2(_156_),
    .ZN(_381_));
 NAND3_X1 _864_ (.A1(_109_),
    .A2(_117_),
    .A3(net60),
    .ZN(_382_));
 NAND2_X2 _865_ (.A1(_381_),
    .A2(_382_),
    .ZN(net51));
 NAND3_X1 _866_ (.A1(_179_),
    .A2(net51),
    .A3(_181_),
    .ZN(_383_));
 OAI21_X1 _867_ (.A(_383_),
    .B1(_183_),
    .B2(net86),
    .ZN(_384_));
 NAND2_X1 _868_ (.A1(_384_),
    .A2(_185_),
    .ZN(_385_));
 AND2_X1 _869_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_386_));
 AOI21_X1 _870_ (.A(_386_),
    .B1(_062_),
    .B2(net17),
    .ZN(_387_));
 NAND2_X1 _871_ (.A1(_385_),
    .A2(_387_),
    .ZN(_018_));
 NAND3_X2 _872_ (.A1(_193_),
    .A2(\dpath.a_lt_b$in1[9] ),
    .A3(_064_),
    .ZN(_388_));
 NAND2_X1 _873_ (.A1(_213_),
    .A2(_214_),
    .ZN(_389_));
 NOR2_X2 _874_ (.A1(_222_),
    .A2(_389_),
    .ZN(_390_));
 NAND3_X2 _875_ (.A1(_390_),
    .A2(_281_),
    .A3(_215_),
    .ZN(_391_));
 INV_X1 _876_ (.A(_286_),
    .ZN(_392_));
 NAND2_X2 _877_ (.A1(_221_),
    .A2(_218_),
    .ZN(_393_));
 NAND2_X1 _878_ (.A1(_393_),
    .A2(_231_),
    .ZN(_394_));
 NAND2_X1 _879_ (.A1(_394_),
    .A2(_281_),
    .ZN(_395_));
 NAND3_X2 _880_ (.A1(_391_),
    .A2(_392_),
    .A3(_395_),
    .ZN(_396_));
 XNOR2_X2 _881_ (.A(_396_),
    .B(_151_),
    .ZN(net52));
 NAND2_X1 _882_ (.A1(net52),
    .A2(_206_),
    .ZN(_397_));
 NAND2_X1 _883_ (.A1(_388_),
    .A2(_397_),
    .ZN(_398_));
 NAND2_X2 _884_ (.A1(_398_),
    .A2(_185_),
    .ZN(_399_));
 AND2_X1 _885_ (.A1(_188_),
    .A2(\dpath.a_lt_b$in0[9] ),
    .ZN(_400_));
 AOI21_X2 _886_ (.A(_400_),
    .B1(_062_),
    .B2(net18),
    .ZN(_401_));
 NAND2_X1 _887_ (.A1(_399_),
    .A2(_401_),
    .ZN(_019_));
 NAND2_X2 _888_ (.A1(_192_),
    .A2(_064_),
    .ZN(_402_));
 BUF_X2 _889_ (.A(_402_),
    .Z(_403_));
 MUX2_X1 _890_ (.A(\dpath.a_lt_b$in0[0] ),
    .B(net1),
    .S(_061_),
    .Z(_404_));
 NAND2_X1 _891_ (.A1(_403_),
    .A2(_404_),
    .ZN(_405_));
 BUF_X2 _892_ (.A(_402_),
    .Z(_406_));
 OAI21_X2 _893_ (.A(_405_),
    .B1(_049_),
    .B2(_406_),
    .ZN(_020_));
 NAND2_X2 _894_ (.A1(_066_),
    .A2(net2),
    .ZN(_407_));
 OAI21_X1 _895_ (.A(_407_),
    .B1(_062_),
    .B2(_143_),
    .ZN(_408_));
 NAND2_X1 _896_ (.A1(_403_),
    .A2(_408_),
    .ZN(_409_));
 OAI21_X1 _897_ (.A(_409_),
    .B1(net73),
    .B2(_406_),
    .ZN(_021_));
 NAND2_X2 _898_ (.A1(_066_),
    .A2(net3),
    .ZN(_410_));
 OAI21_X1 _899_ (.A(_410_),
    .B1(_062_),
    .B2(_139_),
    .ZN(_411_));
 NAND2_X1 _900_ (.A1(_403_),
    .A2(_411_),
    .ZN(_412_));
 OAI21_X2 _901_ (.A(_412_),
    .B1(_036_),
    .B2(_406_),
    .ZN(_022_));
 NAND2_X1 _902_ (.A1(_066_),
    .A2(net4),
    .ZN(_413_));
 BUF_X2 _903_ (.A(_061_),
    .Z(_414_));
 OAI21_X2 _904_ (.A(_413_),
    .B1(_414_),
    .B2(net66),
    .ZN(_415_));
 NAND2_X1 _905_ (.A1(_403_),
    .A2(_415_),
    .ZN(_416_));
 OAI21_X2 _906_ (.A(_416_),
    .B1(net67),
    .B2(_406_),
    .ZN(_023_));
 BUF_X2 _907_ (.A(_402_),
    .Z(_417_));
 NAND2_X1 _908_ (.A1(_066_),
    .A2(net5),
    .ZN(_418_));
 OAI21_X1 _909_ (.A(_418_),
    .B1(_414_),
    .B2(_119_),
    .ZN(_419_));
 NAND2_X1 _910_ (.A1(_417_),
    .A2(_419_),
    .ZN(_420_));
 OAI21_X2 _911_ (.A(_420_),
    .B1(_043_),
    .B2(_406_),
    .ZN(_024_));
 NAND2_X1 _912_ (.A1(_066_),
    .A2(net6),
    .ZN(_421_));
 OAI21_X2 _913_ (.A(_421_),
    .B1(_414_),
    .B2(_131_),
    .ZN(_422_));
 NAND2_X1 _914_ (.A1(_417_),
    .A2(_422_),
    .ZN(_423_));
 OAI21_X1 _915_ (.A(_423_),
    .B1(_042_),
    .B2(_406_),
    .ZN(_025_));
 MUX2_X1 _916_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(net7),
    .S(_061_),
    .Z(_424_));
 NAND2_X2 _917_ (.A1(_417_),
    .A2(_424_),
    .ZN(_425_));
 OAI21_X1 _918_ (.A(_425_),
    .B1(_041_),
    .B2(_406_),
    .ZN(_026_));
 MUX2_X1 _919_ (.A(\dpath.a_lt_b$in0[1] ),
    .B(net12),
    .S(_061_),
    .Z(_426_));
 NAND2_X1 _920_ (.A1(_417_),
    .A2(_426_),
    .ZN(_427_));
 OAI21_X2 _921_ (.A(_427_),
    .B1(_048_),
    .B2(_406_),
    .ZN(_027_));
 NAND2_X2 _922_ (.A1(_066_),
    .A2(net23),
    .ZN(_428_));
 OAI21_X1 _923_ (.A(_428_),
    .B1(_414_),
    .B2(net118),
    .ZN(_429_));
 NAND2_X2 _924_ (.A1(_417_),
    .A2(_429_),
    .ZN(_430_));
 OAI21_X2 _925_ (.A(_430_),
    .B1(_047_),
    .B2(_406_),
    .ZN(_028_));
 NAND2_X1 _926_ (.A1(_066_),
    .A2(net26),
    .ZN(_431_));
 OAI21_X1 _927_ (.A(_431_),
    .B1(_414_),
    .B2(net121),
    .ZN(_432_));
 NAND2_X2 _928_ (.A1(_417_),
    .A2(_432_),
    .ZN(_433_));
 OAI21_X2 _929_ (.A(_433_),
    .B1(_046_),
    .B2(_406_),
    .ZN(_029_));
 NAND2_X1 _930_ (.A1(_066_),
    .A2(net27),
    .ZN(_434_));
 OAI21_X1 _931_ (.A(_434_),
    .B1(_414_),
    .B2(_104_),
    .ZN(_435_));
 NAND2_X1 _932_ (.A1(_417_),
    .A2(_435_),
    .ZN(_436_));
 OAI21_X2 _933_ (.A(_436_),
    .B1(net101),
    .B2(_403_),
    .ZN(_030_));
 NAND2_X2 _934_ (.A1(_061_),
    .A2(net28),
    .ZN(_437_));
 OAI21_X2 _935_ (.A(_437_),
    .B1(_414_),
    .B2(net59),
    .ZN(_438_));
 NAND2_X1 _936_ (.A1(_417_),
    .A2(_438_),
    .ZN(_439_));
 OAI21_X1 _937_ (.A(_439_),
    .B1(net103),
    .B2(_403_),
    .ZN(_031_));
 NAND2_X2 _938_ (.A1(_061_),
    .A2(net29),
    .ZN(_440_));
 OAI21_X1 _939_ (.A(_440_),
    .B1(_414_),
    .B2(net122),
    .ZN(_441_));
 NAND2_X2 _940_ (.A1(_417_),
    .A2(_441_),
    .ZN(_442_));
 OAI21_X1 _941_ (.A(_442_),
    .B1(net123),
    .B2(_403_),
    .ZN(_032_));
 NAND2_X1 _942_ (.A1(_061_),
    .A2(net30),
    .ZN(_443_));
 OAI21_X1 _943_ (.A(_443_),
    .B1(_414_),
    .B2(_090_),
    .ZN(_444_));
 NAND2_X1 _944_ (.A1(_417_),
    .A2(_444_),
    .ZN(_445_));
 OAI21_X1 _945_ (.A(_445_),
    .B1(_051_),
    .B2(_403_),
    .ZN(_033_));
 NAND2_X2 _946_ (.A1(_061_),
    .A2(net31),
    .ZN(_446_));
 OAI21_X1 _947_ (.A(_446_),
    .B1(_414_),
    .B2(net87),
    .ZN(_447_));
 NAND2_X1 _948_ (.A1(_402_),
    .A2(_447_),
    .ZN(_448_));
 OAI21_X1 _949_ (.A(_448_),
    .B1(net85),
    .B2(_403_),
    .ZN(_034_));
 NAND2_X1 _950_ (.A1(_061_),
    .A2(net32),
    .ZN(_449_));
 OAI21_X1 _951_ (.A(_449_),
    .B1(_066_),
    .B2(_149_),
    .ZN(_450_));
 NAND2_X2 _952_ (.A1(_402_),
    .A2(_450_),
    .ZN(_451_));
 OAI21_X1 _953_ (.A(_451_),
    .B1(net88),
    .B2(_403_),
    .ZN(_035_));
 DFF_X1 \ctrl.state.out[0]$_DFF_P_  (.D(_000_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net36),
    .QN(_003_));
 DFF_X1 \ctrl.state.out[1]$_DFF_P_  (.D(_001_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\ctrl.state.out[1] ),
    .QN(_485_));
 DFF_X1 \ctrl.state.out[2]$_DFF_P_  (.D(_002_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\ctrl.state.out[2] ),
    .QN(_484_));
 DFF_X1 \dpath.a_reg.out[0]$_DFFE_PP_  (.D(_004_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[0] ),
    .QN(_483_));
 DFF_X1 \dpath.a_reg.out[10]$_DFFE_PP_  (.D(_005_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[10] ),
    .QN(_482_));
 DFF_X1 \dpath.a_reg.out[11]$_DFFE_PP_  (.D(_006_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[11] ),
    .QN(_481_));
 DFF_X1 \dpath.a_reg.out[12]$_DFFE_PP_  (.D(_007_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[12] ),
    .QN(_480_));
 DFF_X1 \dpath.a_reg.out[13]$_DFFE_PP_  (.D(_008_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[13] ),
    .QN(_479_));
 DFF_X1 \dpath.a_reg.out[14]$_DFFE_PP_  (.D(_009_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[14] ),
    .QN(_478_));
 DFF_X1 \dpath.a_reg.out[15]$_DFFE_PP_  (.D(_010_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[15] ),
    .QN(_477_));
 DFF_X1 \dpath.a_reg.out[1]$_DFFE_PP_  (.D(_011_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[1] ),
    .QN(_476_));
 DFF_X1 \dpath.a_reg.out[2]$_DFFE_PP_  (.D(_012_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[2] ),
    .QN(_475_));
 DFF_X1 \dpath.a_reg.out[3]$_DFFE_PP_  (.D(_013_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in0[3] ),
    .QN(_474_));
 DFF_X1 \dpath.a_reg.out[4]$_DFFE_PP_  (.D(_014_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[4] ),
    .QN(_473_));
 DFF_X1 \dpath.a_reg.out[5]$_DFFE_PP_  (.D(_015_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[5] ),
    .QN(_472_));
 DFF_X1 \dpath.a_reg.out[6]$_DFFE_PP_  (.D(_016_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in0[6] ),
    .QN(_471_));
 DFF_X1 \dpath.a_reg.out[7]$_DFFE_PP_  (.D(_017_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[7] ),
    .QN(_470_));
 DFF_X1 \dpath.a_reg.out[8]$_DFFE_PP_  (.D(_018_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in0[8] ),
    .QN(_469_));
 DFF_X1 \dpath.a_reg.out[9]$_DFFE_PP_  (.D(_019_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in0[9] ),
    .QN(_468_));
 DFF_X1 \dpath.b_reg.out[0]$_DFFE_PP_  (.D(_020_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[0] ),
    .QN(_467_));
 DFF_X1 \dpath.b_reg.out[10]$_DFFE_PP_  (.D(_021_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[10] ),
    .QN(_466_));
 DFF_X1 \dpath.b_reg.out[11]$_DFFE_PP_  (.D(_022_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[11] ),
    .QN(_465_));
 DFF_X1 \dpath.b_reg.out[12]$_DFFE_PP_  (.D(_023_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[12] ),
    .QN(_464_));
 DFF_X1 \dpath.b_reg.out[13]$_DFFE_PP_  (.D(_024_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[13] ),
    .QN(_463_));
 DFF_X1 \dpath.b_reg.out[14]$_DFFE_PP_  (.D(_025_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[14] ),
    .QN(_462_));
 DFF_X1 \dpath.b_reg.out[15]$_DFFE_PP_  (.D(_026_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[15] ),
    .QN(_461_));
 DFF_X1 \dpath.b_reg.out[1]$_DFFE_PP_  (.D(_027_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\dpath.a_lt_b$in1[1] ),
    .QN(_460_));
 DFF_X1 \dpath.b_reg.out[2]$_DFFE_PP_  (.D(_028_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[2] ),
    .QN(_459_));
 DFF_X1 \dpath.b_reg.out[3]$_DFFE_PP_  (.D(_029_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[3] ),
    .QN(_458_));
 DFF_X1 \dpath.b_reg.out[4]$_DFFE_PP_  (.D(_030_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[4] ),
    .QN(_457_));
 DFF_X1 \dpath.b_reg.out[5]$_DFFE_PP_  (.D(_031_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[5] ),
    .QN(_456_));
 DFF_X1 \dpath.b_reg.out[6]$_DFFE_PP_  (.D(_032_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\dpath.a_lt_b$in1[6] ),
    .QN(_455_));
 DFF_X1 \dpath.b_reg.out[7]$_DFFE_PP_  (.D(_033_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[7] ),
    .QN(_454_));
 DFF_X1 \dpath.b_reg.out[8]$_DFFE_PP_  (.D(_034_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\dpath.a_lt_b$in1[8] ),
    .QN(_453_));
 DFF_X1 \dpath.b_reg.out[9]$_DFFE_PP_  (.D(_035_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\dpath.a_lt_b$in1[9] ),
    .QN(_452_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_47 ();
 BUF_X1 input1 (.A(req_msg[0]),
    .Z(net1));
 BUF_X1 input2 (.A(req_msg[10]),
    .Z(net2));
 BUF_X1 input3 (.A(req_msg[11]),
    .Z(net3));
 BUF_X1 input4 (.A(req_msg[12]),
    .Z(net4));
 BUF_X1 input5 (.A(req_msg[13]),
    .Z(net5));
 BUF_X2 input6 (.A(req_msg[14]),
    .Z(net6));
 BUF_X1 input7 (.A(req_msg[15]),
    .Z(net7));
 BUF_X2 input8 (.A(req_msg[16]),
    .Z(net8));
 BUF_X1 input9 (.A(req_msg[17]),
    .Z(net9));
 BUF_X2 input10 (.A(req_msg[18]),
    .Z(net10));
 BUF_X2 input11 (.A(req_msg[19]),
    .Z(net11));
 BUF_X2 input12 (.A(req_msg[1]),
    .Z(net12));
 BUF_X1 input13 (.A(req_msg[20]),
    .Z(net13));
 BUF_X1 input14 (.A(req_msg[21]),
    .Z(net14));
 BUF_X1 input15 (.A(req_msg[22]),
    .Z(net15));
 BUF_X1 input16 (.A(req_msg[23]),
    .Z(net16));
 BUF_X1 input17 (.A(req_msg[24]),
    .Z(net17));
 BUF_X1 input18 (.A(req_msg[25]),
    .Z(net18));
 BUF_X2 input19 (.A(req_msg[26]),
    .Z(net19));
 BUF_X1 input20 (.A(req_msg[27]),
    .Z(net20));
 BUF_X1 input21 (.A(req_msg[28]),
    .Z(net21));
 BUF_X1 input22 (.A(req_msg[29]),
    .Z(net22));
 BUF_X2 input23 (.A(req_msg[2]),
    .Z(net23));
 BUF_X1 input24 (.A(req_msg[30]),
    .Z(net24));
 BUF_X2 input25 (.A(req_msg[31]),
    .Z(net25));
 BUF_X1 input26 (.A(req_msg[3]),
    .Z(net26));
 BUF_X1 input27 (.A(req_msg[4]),
    .Z(net27));
 BUF_X1 input28 (.A(req_msg[5]),
    .Z(net28));
 BUF_X1 input29 (.A(req_msg[6]),
    .Z(net29));
 BUF_X2 input30 (.A(req_msg[7]),
    .Z(net30));
 BUF_X2 input31 (.A(req_msg[8]),
    .Z(net31));
 BUF_X1 input32 (.A(req_msg[9]),
    .Z(net32));
 BUF_X1 input33 (.A(req_val),
    .Z(net33));
 BUF_X1 input34 (.A(reset),
    .Z(net34));
 BUF_X1 input35 (.A(resp_rdy),
    .Z(net35));
 BUF_X1 output36 (.A(net36),
    .Z(req_rdy));
 BUF_X1 output37 (.A(net37),
    .Z(resp_msg[0]));
 BUF_X2 output38 (.A(net38),
    .Z(resp_msg[10]));
 BUF_X1 output39 (.A(net39),
    .Z(resp_msg[11]));
 BUF_X1 output40 (.A(net40),
    .Z(resp_msg[12]));
 BUF_X1 output41 (.A(net41),
    .Z(resp_msg[13]));
 BUF_X1 output42 (.A(net42),
    .Z(resp_msg[14]));
 BUF_X1 output43 (.A(net43),
    .Z(resp_msg[15]));
 BUF_X1 output44 (.A(net44),
    .Z(resp_msg[1]));
 BUF_X1 output45 (.A(net45),
    .Z(resp_msg[2]));
 BUF_X2 output46 (.A(net46),
    .Z(resp_msg[3]));
 BUF_X1 output47 (.A(net47),
    .Z(resp_msg[4]));
 BUF_X1 output48 (.A(net48),
    .Z(resp_msg[5]));
 BUF_X1 output49 (.A(net49),
    .Z(resp_msg[6]));
 BUF_X2 output50 (.A(net50),
    .Z(resp_msg[7]));
 BUF_X1 output51 (.A(net51),
    .Z(resp_msg[8]));
 BUF_X1 output52 (.A(net52),
    .Z(resp_msg[9]));
 BUF_X1 output53 (.A(net53),
    .Z(resp_val));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X2 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X2 clkload0 (.A(clknet_2_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_2_2__leaf_clk));
 INV_X2 clkload2 (.A(clknet_2_3__leaf_clk));
 BUF_X2 rebuffer1 (.A(_128_),
    .Z(net54));
 BUF_X2 rebuffer2 (.A(_128_),
    .Z(net55));
 BUF_X2 rebuffer3 (.A(_226_),
    .Z(net56));
 BUF_X2 rebuffer4 (.A(_101_),
    .Z(net57));
 BUF_X4 rebuffer5 (.A(_234_),
    .Z(net58));
 BUF_X1 rebuffer6 (.A(_100_),
    .Z(net59));
 BUF_X2 rebuffer7 (.A(_157_),
    .Z(net60));
 BUF_X2 rebuffer8 (.A(_223_),
    .Z(net61));
 BUF_X2 rebuffer9 (.A(\dpath.a_lt_b$in0[4] ),
    .Z(net62));
 BUF_X1 rebuffer10 (.A(_083_),
    .Z(net63));
 BUF_X2 rebuffer11 (.A(\dpath.a_lt_b$in0[10] ),
    .Z(net64));
 BUF_X1 rebuffer12 (.A(_221_),
    .Z(net65));
 BUF_X2 rebuffer19 (.A(\dpath.a_lt_b$in0[9] ),
    .Z(net72));
 BUF_X1 rebuffer20 (.A(_037_),
    .Z(net73));
 BUF_X1 rebuffer21 (.A(_144_),
    .Z(net74));
 BUF_X1 rebuffer27 (.A(_159_),
    .Z(net80));
 BUF_X2 rebuffer28 (.A(\dpath.a_lt_b$in0[11] ),
    .Z(net81));
 BUF_X1 rebuffer47 (.A(net69),
    .Z(net100));
 BUF_X1 rebuffer48 (.A(net69),
    .Z(net101));
 BUF_X2 rebuffer49 (.A(_053_),
    .Z(net102));
 BUF_X1 rebuffer50 (.A(_053_),
    .Z(net103));
 BUF_X2 rebuffer61 (.A(_118_),
    .Z(net114));
 BUF_X1 rebuffer62 (.A(_089_),
    .Z(net115));
 BUF_X2 rebuffer63 (.A(_089_),
    .Z(net116));
 BUF_X2 rebuffer64 (.A(\dpath.a_lt_b$in1[2] ),
    .Z(net117));
 BUF_X1 rebuffer66 (.A(\dpath.a_lt_b$in1[3] ),
    .Z(net119));
 BUF_X1 rebuffer67 (.A(_079_),
    .Z(net120));
 BUF_X1 rebuffer68 (.A(_077_),
    .Z(net121));
 BUF_X1 rebuffer69 (.A(_095_),
    .Z(net122));
 BUF_X2 rebuffer70 (.A(_052_),
    .Z(net123));
 BUF_X1 rebuffer71 (.A(net50),
    .Z(net124));
 BUF_X1 rebuffer13 (.A(_125_),
    .Z(net66));
 BUF_X1 rebuffer14 (.A(_044_),
    .Z(net67));
 BUF_X1 rebuffer15 (.A(_044_),
    .Z(net68));
 BUF_X1 rebuffer16 (.A(_054_),
    .Z(net69));
 BUF_X1 rebuffer17 (.A(_106_),
    .Z(net70));
 BUF_X4 rebuffer18 (.A(_199_),
    .Z(net71));
 BUF_X2 rebuffer22 (.A(\dpath.a_lt_b$in0[7] ),
    .Z(net75));
 BUF_X1 rebuffer23 (.A(net38),
    .Z(net76));
 BUF_X2 rebuffer24 (.A(\dpath.a_lt_b$in1[4] ),
    .Z(net77));
 BUF_X1 rebuffer31 (.A(_155_),
    .Z(net84));
 BUF_X1 rebuffer32 (.A(_039_),
    .Z(net85));
 BUF_X1 rebuffer33 (.A(_039_),
    .Z(net86));
 BUF_X1 rebuffer34 (.A(_154_),
    .Z(net87));
 BUF_X1 rebuffer35 (.A(_038_),
    .Z(net88));
 BUF_X1 rebuffer36 (.A(_038_),
    .Z(net89));
 BUF_X1 rebuffer41 (.A(net40),
    .Z(net94));
 BUF_X2 rebuffer44 (.A(_233_),
    .Z(net97));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X4 FILLER_0_17 ();
 FILLCELL_X2 FILLER_0_176 ();
 FILLCELL_X1 FILLER_0_178 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_17 ();
 FILLCELL_X1 FILLER_1_19 ();
 FILLCELL_X1 FILLER_1_54 ();
 FILLCELL_X1 FILLER_1_104 ();
 FILLCELL_X1 FILLER_1_117 ();
 FILLCELL_X1 FILLER_1_146 ();
 FILLCELL_X8 FILLER_1_169 ();
 FILLCELL_X2 FILLER_1_177 ();
 FILLCELL_X2 FILLER_2_1 ();
 FILLCELL_X1 FILLER_2_3 ();
 FILLCELL_X4 FILLER_2_21 ();
 FILLCELL_X2 FILLER_2_25 ();
 FILLCELL_X1 FILLER_2_38 ();
 FILLCELL_X1 FILLER_2_42 ();
 FILLCELL_X1 FILLER_2_69 ();
 FILLCELL_X8 FILLER_2_167 ();
 FILLCELL_X4 FILLER_2_175 ();
 FILLCELL_X8 FILLER_3_1 ();
 FILLCELL_X1 FILLER_3_9 ();
 FILLCELL_X4 FILLER_3_17 ();
 FILLCELL_X8 FILLER_3_25 ();
 FILLCELL_X2 FILLER_3_33 ();
 FILLCELL_X1 FILLER_3_35 ();
 FILLCELL_X4 FILLER_3_40 ();
 FILLCELL_X2 FILLER_3_67 ();
 FILLCELL_X1 FILLER_3_108 ();
 FILLCELL_X2 FILLER_3_168 ();
 FILLCELL_X2 FILLER_3_176 ();
 FILLCELL_X1 FILLER_3_178 ();
 FILLCELL_X16 FILLER_4_4 ();
 FILLCELL_X8 FILLER_4_20 ();
 FILLCELL_X2 FILLER_4_32 ();
 FILLCELL_X2 FILLER_4_45 ();
 FILLCELL_X2 FILLER_4_75 ();
 FILLCELL_X2 FILLER_4_84 ();
 FILLCELL_X1 FILLER_4_131 ();
 FILLCELL_X1 FILLER_4_178 ();
 FILLCELL_X16 FILLER_5_1 ();
 FILLCELL_X2 FILLER_5_37 ();
 FILLCELL_X1 FILLER_5_39 ();
 FILLCELL_X2 FILLER_5_47 ();
 FILLCELL_X1 FILLER_5_49 ();
 FILLCELL_X4 FILLER_5_61 ();
 FILLCELL_X1 FILLER_5_65 ();
 FILLCELL_X1 FILLER_5_97 ();
 FILLCELL_X1 FILLER_5_102 ();
 FILLCELL_X4 FILLER_5_173 ();
 FILLCELL_X2 FILLER_5_177 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X4 FILLER_6_9 ();
 FILLCELL_X2 FILLER_6_16 ();
 FILLCELL_X1 FILLER_6_18 ();
 FILLCELL_X8 FILLER_6_22 ();
 FILLCELL_X4 FILLER_6_30 ();
 FILLCELL_X2 FILLER_6_34 ();
 FILLCELL_X1 FILLER_6_49 ();
 FILLCELL_X4 FILLER_6_55 ();
 FILLCELL_X2 FILLER_6_66 ();
 FILLCELL_X8 FILLER_6_72 ();
 FILLCELL_X4 FILLER_6_80 ();
 FILLCELL_X1 FILLER_6_84 ();
 FILLCELL_X1 FILLER_6_88 ();
 FILLCELL_X2 FILLER_6_93 ();
 FILLCELL_X1 FILLER_6_99 ();
 FILLCELL_X1 FILLER_6_160 ();
 FILLCELL_X2 FILLER_6_177 ();
 FILLCELL_X4 FILLER_7_10 ();
 FILLCELL_X1 FILLER_7_14 ();
 FILLCELL_X8 FILLER_7_32 ();
 FILLCELL_X4 FILLER_7_40 ();
 FILLCELL_X1 FILLER_7_44 ();
 FILLCELL_X2 FILLER_7_52 ();
 FILLCELL_X1 FILLER_7_54 ();
 FILLCELL_X4 FILLER_7_78 ();
 FILLCELL_X2 FILLER_7_82 ();
 FILLCELL_X1 FILLER_7_84 ();
 FILLCELL_X1 FILLER_7_99 ();
 FILLCELL_X2 FILLER_7_105 ();
 FILLCELL_X8 FILLER_8_23 ();
 FILLCELL_X2 FILLER_8_38 ();
 FILLCELL_X1 FILLER_8_40 ();
 FILLCELL_X8 FILLER_8_58 ();
 FILLCELL_X8 FILLER_8_71 ();
 FILLCELL_X1 FILLER_8_79 ();
 FILLCELL_X2 FILLER_8_83 ();
 FILLCELL_X1 FILLER_8_89 ();
 FILLCELL_X2 FILLER_8_110 ();
 FILLCELL_X2 FILLER_9_1 ();
 FILLCELL_X2 FILLER_9_11 ();
 FILLCELL_X1 FILLER_9_18 ();
 FILLCELL_X2 FILLER_9_23 ();
 FILLCELL_X8 FILLER_9_28 ();
 FILLCELL_X2 FILLER_9_39 ();
 FILLCELL_X1 FILLER_9_41 ();
 FILLCELL_X8 FILLER_9_50 ();
 FILLCELL_X4 FILLER_9_58 ();
 FILLCELL_X2 FILLER_9_62 ();
 FILLCELL_X4 FILLER_9_71 ();
 FILLCELL_X2 FILLER_9_75 ();
 FILLCELL_X1 FILLER_9_77 ();
 FILLCELL_X2 FILLER_9_82 ();
 FILLCELL_X2 FILLER_9_168 ();
 FILLCELL_X1 FILLER_9_178 ();
 FILLCELL_X2 FILLER_10_7 ();
 FILLCELL_X2 FILLER_10_15 ();
 FILLCELL_X4 FILLER_10_29 ();
 FILLCELL_X2 FILLER_10_33 ();
 FILLCELL_X4 FILLER_10_58 ();
 FILLCELL_X4 FILLER_10_80 ();
 FILLCELL_X2 FILLER_10_84 ();
 FILLCELL_X4 FILLER_10_89 ();
 FILLCELL_X1 FILLER_10_93 ();
 FILLCELL_X2 FILLER_11_1 ();
 FILLCELL_X1 FILLER_11_3 ();
 FILLCELL_X2 FILLER_11_21 ();
 FILLCELL_X1 FILLER_11_23 ();
 FILLCELL_X4 FILLER_11_31 ();
 FILLCELL_X2 FILLER_11_35 ();
 FILLCELL_X1 FILLER_11_37 ();
 FILLCELL_X8 FILLER_11_43 ();
 FILLCELL_X4 FILLER_11_61 ();
 FILLCELL_X1 FILLER_11_78 ();
 FILLCELL_X8 FILLER_11_92 ();
 FILLCELL_X1 FILLER_11_142 ();
 FILLCELL_X2 FILLER_11_177 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X8 FILLER_12_17 ();
 FILLCELL_X2 FILLER_12_25 ();
 FILLCELL_X1 FILLER_12_27 ();
 FILLCELL_X2 FILLER_12_49 ();
 FILLCELL_X2 FILLER_12_70 ();
 FILLCELL_X4 FILLER_12_95 ();
 FILLCELL_X1 FILLER_12_99 ();
 FILLCELL_X2 FILLER_12_177 ();
 FILLCELL_X8 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_9 ();
 FILLCELL_X4 FILLER_13_33 ();
 FILLCELL_X1 FILLER_13_37 ();
 FILLCELL_X1 FILLER_13_52 ();
 FILLCELL_X2 FILLER_13_68 ();
 FILLCELL_X1 FILLER_13_77 ();
 FILLCELL_X1 FILLER_13_88 ();
 FILLCELL_X1 FILLER_13_93 ();
 FILLCELL_X1 FILLER_13_142 ();
 FILLCELL_X1 FILLER_13_174 ();
 FILLCELL_X1 FILLER_13_178 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X4 FILLER_14_9 ();
 FILLCELL_X4 FILLER_14_16 ();
 FILLCELL_X1 FILLER_14_20 ();
 FILLCELL_X2 FILLER_14_53 ();
 FILLCELL_X1 FILLER_14_58 ();
 FILLCELL_X1 FILLER_14_62 ();
 FILLCELL_X1 FILLER_14_81 ();
 FILLCELL_X1 FILLER_14_89 ();
 FILLCELL_X2 FILLER_14_95 ();
 FILLCELL_X1 FILLER_14_109 ();
 FILLCELL_X8 FILLER_14_169 ();
 FILLCELL_X2 FILLER_14_177 ();
 FILLCELL_X1 FILLER_15_4 ();
 FILLCELL_X1 FILLER_15_26 ();
 FILLCELL_X2 FILLER_15_30 ();
 FILLCELL_X1 FILLER_15_112 ();
 FILLCELL_X16 FILLER_15_159 ();
 FILLCELL_X4 FILLER_15_175 ();
 FILLCELL_X4 FILLER_16_1 ();
 FILLCELL_X1 FILLER_16_5 ();
 FILLCELL_X8 FILLER_16_9 ();
 FILLCELL_X4 FILLER_16_17 ();
 FILLCELL_X2 FILLER_16_21 ();
 FILLCELL_X1 FILLER_16_48 ();
 FILLCELL_X2 FILLER_16_69 ();
 FILLCELL_X2 FILLER_16_74 ();
 FILLCELL_X1 FILLER_16_80 ();
 FILLCELL_X1 FILLER_16_107 ();
 FILLCELL_X16 FILLER_16_155 ();
 FILLCELL_X8 FILLER_16_171 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_5 ();
 FILLCELL_X1 FILLER_17_7 ();
 FILLCELL_X16 FILLER_17_11 ();
 FILLCELL_X4 FILLER_17_27 ();
 FILLCELL_X1 FILLER_17_31 ();
 FILLCELL_X2 FILLER_17_35 ();
 FILLCELL_X1 FILLER_17_50 ();
 FILLCELL_X2 FILLER_17_60 ();
 FILLCELL_X2 FILLER_17_79 ();
 FILLCELL_X1 FILLER_17_81 ();
 FILLCELL_X1 FILLER_17_111 ();
 FILLCELL_X16 FILLER_17_159 ();
 FILLCELL_X4 FILLER_17_175 ();
 FILLCELL_X16 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_17 ();
 FILLCELL_X2 FILLER_18_21 ();
 FILLCELL_X16 FILLER_18_26 ();
 FILLCELL_X2 FILLER_18_45 ();
 FILLCELL_X1 FILLER_18_47 ();
 FILLCELL_X1 FILLER_18_83 ();
 FILLCELL_X4 FILLER_18_87 ();
 FILLCELL_X2 FILLER_18_91 ();
 FILLCELL_X1 FILLER_18_93 ();
 FILLCELL_X1 FILLER_18_148 ();
 FILLCELL_X16 FILLER_18_157 ();
 FILLCELL_X4 FILLER_18_173 ();
 FILLCELL_X2 FILLER_18_177 ();
 FILLCELL_X16 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_17 ();
 FILLCELL_X1 FILLER_19_21 ();
 FILLCELL_X2 FILLER_19_26 ();
 FILLCELL_X1 FILLER_19_28 ();
 FILLCELL_X2 FILLER_19_57 ();
 FILLCELL_X1 FILLER_19_59 ();
 FILLCELL_X2 FILLER_19_86 ();
 FILLCELL_X1 FILLER_19_88 ();
 FILLCELL_X4 FILLER_19_92 ();
 FILLCELL_X2 FILLER_19_96 ();
 FILLCELL_X1 FILLER_19_109 ();
 FILLCELL_X1 FILLER_19_113 ();
 FILLCELL_X1 FILLER_19_124 ();
 FILLCELL_X1 FILLER_19_140 ();
 FILLCELL_X16 FILLER_19_151 ();
 FILLCELL_X8 FILLER_19_167 ();
 FILLCELL_X4 FILLER_19_175 ();
 FILLCELL_X2 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_6 ();
 FILLCELL_X1 FILLER_20_8 ();
 FILLCELL_X4 FILLER_20_33 ();
 FILLCELL_X2 FILLER_20_37 ();
 FILLCELL_X2 FILLER_20_51 ();
 FILLCELL_X1 FILLER_20_94 ();
 FILLCELL_X1 FILLER_20_123 ();
 FILLCELL_X2 FILLER_20_136 ();
 FILLCELL_X32 FILLER_20_144 ();
 FILLCELL_X2 FILLER_20_176 ();
 FILLCELL_X1 FILLER_20_178 ();
 FILLCELL_X16 FILLER_21_1 ();
 FILLCELL_X8 FILLER_21_17 ();
 FILLCELL_X2 FILLER_21_25 ();
 FILLCELL_X4 FILLER_21_34 ();
 FILLCELL_X2 FILLER_21_38 ();
 FILLCELL_X1 FILLER_21_40 ();
 FILLCELL_X8 FILLER_21_48 ();
 FILLCELL_X1 FILLER_21_56 ();
 FILLCELL_X1 FILLER_21_63 ();
 FILLCELL_X1 FILLER_21_72 ();
 FILLCELL_X4 FILLER_21_87 ();
 FILLCELL_X2 FILLER_21_91 ();
 FILLCELL_X2 FILLER_21_116 ();
 FILLCELL_X32 FILLER_21_145 ();
 FILLCELL_X2 FILLER_21_177 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X2 FILLER_22_17 ();
 FILLCELL_X1 FILLER_22_19 ();
 FILLCELL_X2 FILLER_22_54 ();
 FILLCELL_X2 FILLER_22_75 ();
 FILLCELL_X1 FILLER_22_77 ();
 FILLCELL_X8 FILLER_22_105 ();
 FILLCELL_X4 FILLER_22_113 ();
 FILLCELL_X2 FILLER_22_117 ();
 FILLCELL_X1 FILLER_22_119 ();
 FILLCELL_X32 FILLER_22_136 ();
 FILLCELL_X8 FILLER_22_168 ();
 FILLCELL_X2 FILLER_22_176 ();
 FILLCELL_X1 FILLER_22_178 ();
 FILLCELL_X16 FILLER_23_1 ();
 FILLCELL_X4 FILLER_23_17 ();
 FILLCELL_X2 FILLER_23_21 ();
 FILLCELL_X1 FILLER_23_23 ();
 FILLCELL_X4 FILLER_23_31 ();
 FILLCELL_X1 FILLER_23_35 ();
 FILLCELL_X8 FILLER_23_52 ();
 FILLCELL_X2 FILLER_23_60 ();
 FILLCELL_X4 FILLER_23_75 ();
 FILLCELL_X4 FILLER_23_82 ();
 FILLCELL_X4 FILLER_23_92 ();
 FILLCELL_X2 FILLER_23_96 ();
 FILLCELL_X1 FILLER_23_98 ();
 FILLCELL_X2 FILLER_23_102 ();
 FILLCELL_X8 FILLER_23_110 ();
 FILLCELL_X2 FILLER_23_121 ();
 FILLCELL_X1 FILLER_23_123 ();
 FILLCELL_X32 FILLER_23_127 ();
 FILLCELL_X16 FILLER_23_159 ();
 FILLCELL_X4 FILLER_23_175 ();
endmodule
